module PUFMux256(i_D, i_Sel, o_Q);

    input [255:0] i_D;
    input [7:0] i_Sel;
    output reg o_Q;

    always@(*) begin
        case(i_Sel)
            8'b00000000: o_Q <= i_D[0];
            8'b00000001: o_Q <= i_D[1];
            8'b00000010: o_Q <= i_D[2];
            8'b00000011: o_Q <= i_D[3];
            8'b00000100: o_Q <= i_D[4];
            8'b00000101: o_Q <= i_D[5];
            8'b00000110: o_Q <= i_D[6];
            8'b00000111: o_Q <= i_D[7];
            8'b00001000: o_Q <= i_D[8];
            8'b00001001: o_Q <= i_D[9];
            8'b00001010: o_Q <= i_D[10];
            8'b00001011: o_Q <= i_D[11];
            8'b00001100: o_Q <= i_D[12];
            8'b00001101: o_Q <= i_D[13];
            8'b00001110: o_Q <= i_D[14];
            8'b00001111: o_Q <= i_D[15];
            8'b00010000: o_Q <= i_D[16];
            8'b00010001: o_Q <= i_D[17];
            8'b00010010: o_Q <= i_D[18];
            8'b00010011: o_Q <= i_D[19];
            8'b00010100: o_Q <= i_D[20];
            8'b00010101: o_Q <= i_D[21];
            8'b00010110: o_Q <= i_D[22];
            8'b00010111: o_Q <= i_D[23];
            8'b00011000: o_Q <= i_D[24];
            8'b00011001: o_Q <= i_D[25];
            8'b00011010: o_Q <= i_D[26];
            8'b00011011: o_Q <= i_D[27];
            8'b00011100: o_Q <= i_D[28];
            8'b00011101: o_Q <= i_D[29];
            8'b00011110: o_Q <= i_D[30];
            8'b00011111: o_Q <= i_D[31];
            8'b00100000: o_Q <= i_D[32];
            8'b00100001: o_Q <= i_D[33];
            8'b00100010: o_Q <= i_D[34];
            8'b00100011: o_Q <= i_D[35];
            8'b00100100: o_Q <= i_D[36];
            8'b00100101: o_Q <= i_D[37];
            8'b00100110: o_Q <= i_D[38];
            8'b00100111: o_Q <= i_D[39];
            8'b00101000: o_Q <= i_D[40];
            8'b00101001: o_Q <= i_D[41];
            8'b00101010: o_Q <= i_D[42];
            8'b00101011: o_Q <= i_D[43];
            8'b00101100: o_Q <= i_D[44];
            8'b00101101: o_Q <= i_D[45];
            8'b00101110: o_Q <= i_D[46];
            8'b00101111: o_Q <= i_D[47];
            8'b00110000: o_Q <= i_D[48];
            8'b00110001: o_Q <= i_D[49];
            8'b00110010: o_Q <= i_D[50];
            8'b00110011: o_Q <= i_D[51];
            8'b00110100: o_Q <= i_D[52];
            8'b00110101: o_Q <= i_D[53];
            8'b00110110: o_Q <= i_D[54];
            8'b00110111: o_Q <= i_D[55];
            8'b00111000: o_Q <= i_D[56];
            8'b00111001: o_Q <= i_D[57];
            8'b00111010: o_Q <= i_D[58];
            8'b00111011: o_Q <= i_D[59];
            8'b00111100: o_Q <= i_D[60];
            8'b00111101: o_Q <= i_D[61];
            8'b00111110: o_Q <= i_D[62];
            8'b00111111: o_Q <= i_D[63];
            8'b01000000: o_Q <= i_D[64];
            8'b01000001: o_Q <= i_D[65];
            8'b01000010: o_Q <= i_D[66];
            8'b01000011: o_Q <= i_D[67];
            8'b01000100: o_Q <= i_D[68];
            8'b01000101: o_Q <= i_D[69];
            8'b01000110: o_Q <= i_D[70];
            8'b01000111: o_Q <= i_D[71];
            8'b01001000: o_Q <= i_D[72];
            8'b01001001: o_Q <= i_D[73];
            8'b01001010: o_Q <= i_D[74];
            8'b01001011: o_Q <= i_D[75];
            8'b01001100: o_Q <= i_D[76];
            8'b01001101: o_Q <= i_D[77];
            8'b01001110: o_Q <= i_D[78];
            8'b01001111: o_Q <= i_D[79];
            8'b01010000: o_Q <= i_D[80];
            8'b01010001: o_Q <= i_D[81];
            8'b01010010: o_Q <= i_D[82];
            8'b01010011: o_Q <= i_D[83];
            8'b01010100: o_Q <= i_D[84];
            8'b01010101: o_Q <= i_D[85];
            8'b01010110: o_Q <= i_D[86];
            8'b01010111: o_Q <= i_D[87];
            8'b01011000: o_Q <= i_D[88];
            8'b01011001: o_Q <= i_D[89];
            8'b01011010: o_Q <= i_D[90];
            8'b01011011: o_Q <= i_D[91];
            8'b01011100: o_Q <= i_D[92];
            8'b01011101: o_Q <= i_D[93];
            8'b01011110: o_Q <= i_D[94];
            8'b01011111: o_Q <= i_D[95];
            8'b01100000: o_Q <= i_D[96];
            8'b01100001: o_Q <= i_D[97];
            8'b01100010: o_Q <= i_D[98];
            8'b01100011: o_Q <= i_D[99];
            8'b01100100: o_Q <= i_D[100];
            8'b01100101: o_Q <= i_D[101];
            8'b01100110: o_Q <= i_D[102];
            8'b01100111: o_Q <= i_D[103];
            8'b01101000: o_Q <= i_D[104];
            8'b01101001: o_Q <= i_D[105];
            8'b01101010: o_Q <= i_D[106];
            8'b01101011: o_Q <= i_D[107];
            8'b01101100: o_Q <= i_D[108];
            8'b01101101: o_Q <= i_D[109];
            8'b01101110: o_Q <= i_D[110];
            8'b01101111: o_Q <= i_D[111];
            8'b01110000: o_Q <= i_D[112];
            8'b01110001: o_Q <= i_D[113];
            8'b01110010: o_Q <= i_D[114];
            8'b01110011: o_Q <= i_D[115];
            8'b01110100: o_Q <= i_D[116];
            8'b01110101: o_Q <= i_D[117];
            8'b01110110: o_Q <= i_D[118];
            8'b01110111: o_Q <= i_D[119];
            8'b01111000: o_Q <= i_D[120];
            8'b01111001: o_Q <= i_D[121];
            8'b01111010: o_Q <= i_D[122];
            8'b01111011: o_Q <= i_D[123];
            8'b01111100: o_Q <= i_D[124];
            8'b01111101: o_Q <= i_D[125];
            8'b01111110: o_Q <= i_D[126];
            8'b01111111: o_Q <= i_D[127];
            8'b10000000: o_Q <= i_D[128];
            8'b10000001: o_Q <= i_D[129];
            8'b10000010: o_Q <= i_D[130];
            8'b10000011: o_Q <= i_D[131];
            8'b10000100: o_Q <= i_D[132];
            8'b10000101: o_Q <= i_D[133];
            8'b10000110: o_Q <= i_D[134];
            8'b10000111: o_Q <= i_D[135];
            8'b10001000: o_Q <= i_D[136];
            8'b10001001: o_Q <= i_D[137];
            8'b10001010: o_Q <= i_D[138];
            8'b10001011: o_Q <= i_D[139];
            8'b10001100: o_Q <= i_D[140];
            8'b10001101: o_Q <= i_D[141];
            8'b10001110: o_Q <= i_D[142];
            8'b10001111: o_Q <= i_D[143];
            8'b10010000: o_Q <= i_D[144];
            8'b10010001: o_Q <= i_D[145];
            8'b10010010: o_Q <= i_D[146];
            8'b10010011: o_Q <= i_D[147];
            8'b10010100: o_Q <= i_D[148];
            8'b10010101: o_Q <= i_D[149];
            8'b10010110: o_Q <= i_D[150];
            8'b10010111: o_Q <= i_D[151];
            8'b10011000: o_Q <= i_D[152];
            8'b10011001: o_Q <= i_D[153];
            8'b10011010: o_Q <= i_D[154];
            8'b10011011: o_Q <= i_D[155];
            8'b10011100: o_Q <= i_D[156];
            8'b10011101: o_Q <= i_D[157];
            8'b10011110: o_Q <= i_D[158];
            8'b10011111: o_Q <= i_D[159];
            8'b10100000: o_Q <= i_D[160];
            8'b10100001: o_Q <= i_D[161];
            8'b10100010: o_Q <= i_D[162];
            8'b10100011: o_Q <= i_D[163];
            8'b10100100: o_Q <= i_D[164];
            8'b10100101: o_Q <= i_D[165];
            8'b10100110: o_Q <= i_D[166];
            8'b10100111: o_Q <= i_D[167];
            8'b10101000: o_Q <= i_D[168];
            8'b10101001: o_Q <= i_D[169];
            8'b10101010: o_Q <= i_D[170];
            8'b10101011: o_Q <= i_D[171];
            8'b10101100: o_Q <= i_D[172];
            8'b10101101: o_Q <= i_D[173];
            8'b10101110: o_Q <= i_D[174];
            8'b10101111: o_Q <= i_D[175];
            8'b10110000: o_Q <= i_D[176];
            8'b10110001: o_Q <= i_D[177];
            8'b10110010: o_Q <= i_D[178];
            8'b10110011: o_Q <= i_D[179];
            8'b10110100: o_Q <= i_D[180];
            8'b10110101: o_Q <= i_D[181];
            8'b10110110: o_Q <= i_D[182];
            8'b10110111: o_Q <= i_D[183];
            8'b10111000: o_Q <= i_D[184];
            8'b10111001: o_Q <= i_D[185];
            8'b10111010: o_Q <= i_D[186];
            8'b10111011: o_Q <= i_D[187];
            8'b10111100: o_Q <= i_D[188];
            8'b10111101: o_Q <= i_D[189];
            8'b10111110: o_Q <= i_D[190];
            8'b10111111: o_Q <= i_D[191];
            8'b11000000: o_Q <= i_D[192];
            8'b11000001: o_Q <= i_D[193];
            8'b11000010: o_Q <= i_D[194];
            8'b11000011: o_Q <= i_D[195];
            8'b11000100: o_Q <= i_D[196];
            8'b11000101: o_Q <= i_D[197];
            8'b11000110: o_Q <= i_D[198];
            8'b11000111: o_Q <= i_D[199];
            8'b11001000: o_Q <= i_D[200];
            8'b11001001: o_Q <= i_D[201];
            8'b11001010: o_Q <= i_D[202];
            8'b11001011: o_Q <= i_D[203];
            8'b11001100: o_Q <= i_D[204];
            8'b11001101: o_Q <= i_D[205];
            8'b11001110: o_Q <= i_D[206];
            8'b11001111: o_Q <= i_D[207];
            8'b11010000: o_Q <= i_D[208];
            8'b11010001: o_Q <= i_D[209];
            8'b11010010: o_Q <= i_D[210];
            8'b11010011: o_Q <= i_D[211];
            8'b11010100: o_Q <= i_D[212];
            8'b11010101: o_Q <= i_D[213];
            8'b11010110: o_Q <= i_D[214];
            8'b11010111: o_Q <= i_D[215];
            8'b11011000: o_Q <= i_D[216];
            8'b11011001: o_Q <= i_D[217];
            8'b11011010: o_Q <= i_D[218];
            8'b11011011: o_Q <= i_D[219];
            8'b11011100: o_Q <= i_D[220];
            8'b11011101: o_Q <= i_D[221];
            8'b11011110: o_Q <= i_D[222];
            8'b11011111: o_Q <= i_D[223];
            8'b11100000: o_Q <= i_D[224];
            8'b11100001: o_Q <= i_D[225];
            8'b11100010: o_Q <= i_D[226];
            8'b11100011: o_Q <= i_D[227];
            8'b11100100: o_Q <= i_D[228];
            8'b11100101: o_Q <= i_D[229];
            8'b11100110: o_Q <= i_D[230];
            8'b11100111: o_Q <= i_D[231];
            8'b11101000: o_Q <= i_D[232];
            8'b11101001: o_Q <= i_D[233];
            8'b11101010: o_Q <= i_D[234];
            8'b11101011: o_Q <= i_D[235];
            8'b11101100: o_Q <= i_D[236];
            8'b11101101: o_Q <= i_D[237];
            8'b11101110: o_Q <= i_D[238];
            8'b11101111: o_Q <= i_D[239];
            8'b11110000: o_Q <= i_D[240];
            8'b11110001: o_Q <= i_D[241];
            8'b11110010: o_Q <= i_D[242];
            8'b11110011: o_Q <= i_D[243];
            8'b11110100: o_Q <= i_D[244];
            8'b11110101: o_Q <= i_D[245];
            8'b11110110: o_Q <= i_D[246];
            8'b11110111: o_Q <= i_D[247];
            8'b11111000: o_Q <= i_D[248];
            8'b11111001: o_Q <= i_D[249];
            8'b11111010: o_Q <= i_D[250];
            8'b11111011: o_Q <= i_D[251];
            8'b11111100: o_Q <= i_D[252];
            8'b11111101: o_Q <= i_D[253];
            8'b11111110: o_Q <= i_D[254];
            8'b11111111: o_Q <= i_D[255];
            default: o_Q <= i_D[255];

        endcase
    end

endmodule
